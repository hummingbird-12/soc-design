* SPICE3 file created from s161577NOT.ext - technology: scmos

.option scale=1u
.include scmos_spice.prm

M1000 F A Vdd Vdd pfet w=11 l=2
+  ad=55 pd=32 as=55 ps=32
M1001 F A Gnd Gnd nfet w=11 l=2
+  ad=55 pd=32 as=55 ps=32

V11 Vdd Gnd 3.3
V01 A Gnd PULSE(0 3.3 1ns 0.2ns 0.2ns 4ns 8.2ns)

.TRAN 0.1ns 10ns

.end
