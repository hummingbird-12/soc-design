magic
tech scmos
timestamp 1601668355
<< polysilicon >>
rect -6 14 -4 16
rect -6 0 -4 10
rect -6 -6 -4 -4
<< ndiffusion >>
rect -7 -4 -6 0
rect -4 -4 -3 0
<< pdiffusion >>
rect -7 10 -6 14
rect -4 10 -3 14
<< metal1 >>
rect -11 14 -7 16
rect -3 0 1 10
rect -11 -6 -7 -4
<< ntransistor >>
rect -6 -4 -4 0
<< ptransistor >>
rect -6 10 -4 14
<< ndcontact >>
rect -11 -4 -7 0
rect -3 -4 1 0
<< pdcontact >>
rect -11 10 -7 14
rect -3 10 1 14
<< psubstratepcontact >>
rect -15 -4 -11 0
<< nsubstratencontact >>
rect -15 10 -11 14
<< labels >>
rlabel polysilicon -5 8 -5 8 1 A
rlabel metal1 -9 15 -9 15 5 Vdd!
rlabel metal1 -9 -5 -9 -5 1 Gnd!
rlabel metal1 -1 8 -1 8 7 F
<< end >>
