* SPICE3 file created from s161577NAND2.ext - technology: scmos

.option scale=1u
.include scmos_spice.prm

M1000 F A Vdd Vdd pfet w=27 l=2
+  ad=162 pd=66 as=270 ps=128
M1001 Vdd B F Vdd pfet w=27 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_n6_n15# A Gnd Gnd nfet w=11 l=2
+  ad=66 pd=34 as=55 ps=32
M1003 F B a_n6_n15# Gnd nfet w=11 l=2
+  ad=55 pd=32 as=0 ps=0

V11 Vdd Gnd 3.3
* V01 A Gnd PULSE(0 3.3 1ns 0.2ns 0.2ns 8ns 16.2ns)
* V02 B Gnd PULSE(0 3.3 5ns 0.2ns 0.2ns 8ns 16.2ns)
V01 A Gnd EXP(0 3.3 4ns 0.2ns 16ns 0.2ns)
V02 B Gnd EXP(0 3.3 10ns 0.2ns 22ns 0.2ns)

.TRAN 0.1ns 25ns

.end
