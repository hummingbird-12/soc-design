magic
tech scmos
timestamp 1601658634
<< polysilicon >>
rect 3 -6 5 -4
rect 11 -6 13 -4
<< metal1 >>
rect -18 3 2 7
rect -26 -7 -22 -3
rect -15 -4 10 0
rect -18 -11 2 -7
<< metal2 >>
rect -19 -4 -15 0
<< polycontact >>
rect -19 -4 -15 0
use s161577NOT_44-25  s161577NOT_44-25_0
timestamp 1601633939
transform 1 0 56 0 1 -2
box -82 -11 -66 11
use s161577NOR_44-25  s161577NOR_44-25_0
timestamp 1601643379
transform 1 0 10 0 1 0
box -16 -16 8 9
<< labels >>
rlabel polysilicon 4 -5 4 -5 1 A
rlabel polysilicon 12 -5 12 -5 1 B
rlabel metal1 -24 -5 -24 -5 3 F
rlabel metal1 -8 -9 -8 -9 1 Gnd!
rlabel metal1 -8 5 -8 5 5 Vdd!
rlabel metal1 8 -2 8 -2 1 NOT_F
<< end >>
