magic
tech scmos
timestamp 1601495434
<< polysilicon >>
rect -8 17 -6 19
rect 0 17 2 19
rect -8 -4 -6 6
rect 0 -4 2 6
rect -8 -17 -6 -15
rect 0 -17 2 -15
<< ndiffusion >>
rect -13 -11 -8 -4
rect -9 -15 -8 -11
rect -6 -15 0 -4
rect 2 -8 3 -4
rect 2 -15 7 -8
<< pdiffusion >>
rect -9 13 -8 17
rect -13 6 -8 13
rect -6 10 0 17
rect -6 6 -5 10
rect -1 6 0 10
rect 2 13 3 17
rect 2 6 7 13
<< metal1 >>
rect -9 13 3 17
rect 7 13 10 17
rect -4 -4 -1 6
rect -4 -7 3 -4
rect -9 -15 10 -11
<< ntransistor >>
rect -8 -15 -6 -4
rect 0 -15 2 -4
<< ptransistor >>
rect -8 6 -6 17
rect 0 6 2 17
<< ndcontact >>
rect -13 -15 -9 -11
rect 3 -8 7 -4
<< pdcontact >>
rect -13 13 -9 17
rect -5 6 -1 10
rect 3 13 7 17
<< psubstratepcontact >>
rect -17 -15 -13 -11
<< nsubstratencontact >>
rect -17 13 -13 17
<< labels >>
rlabel metal1 8 15 8 15 6 Vdd!
rlabel metal1 8 -13 8 -13 7 Gnd!
rlabel polysilicon -7 2 -7 2 1 A
rlabel polysilicon 1 2 1 2 1 B
rlabel metal1 -2 2 -2 2 1 F
<< end >>
