magic
tech scmos
timestamp 1601497156
<< polysilicon >>
rect -1 28 1 30
rect -1 -9 1 1
rect -1 -22 1 -20
<< ndiffusion >>
rect -6 -16 -1 -9
rect -2 -20 -1 -16
rect 1 -13 2 -9
rect 1 -20 6 -13
<< pdiffusion >>
rect -2 24 -1 28
rect -6 1 -1 24
rect 1 5 6 28
rect 1 1 2 5
<< metal1 >>
rect -2 24 9 28
rect 3 -9 6 1
rect -2 -20 9 -16
<< ntransistor >>
rect -1 -20 1 -9
<< ptransistor >>
rect -1 1 1 28
<< ndcontact >>
rect -6 -20 -2 -16
rect 2 -13 6 -9
<< pdcontact >>
rect -6 24 -2 28
rect 2 1 6 5
<< psubstratepcontact >>
rect -10 -20 -6 -16
<< nsubstratencontact >>
rect -10 24 -6 28
<< labels >>
rlabel metal1 7 -18 7 -18 7 Gnd!
rlabel polysilicon 0 -2 0 -2 1 A
rlabel metal1 5 -2 5 -2 7 F
rlabel metal1 7 26 7 26 6 Vdd!
<< end >>
