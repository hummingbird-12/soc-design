magic
tech scmos
timestamp 1601458543
<< polysilicon >>
rect -1 12 1 14
rect -1 -9 1 1
rect -1 -22 1 -20
<< ndiffusion >>
rect -6 -16 -1 -9
rect -2 -20 -1 -16
rect 1 -13 2 -9
rect 1 -20 6 -13
<< pdiffusion >>
rect -2 8 -1 12
rect -6 1 -1 8
rect 1 5 6 12
rect 1 1 2 5
<< metal1 >>
rect -2 8 9 12
rect 3 -9 6 1
rect -2 -20 9 -16
<< ntransistor >>
rect -1 -20 1 -9
<< ptransistor >>
rect -1 1 1 12
<< ndcontact >>
rect -6 -20 -2 -16
rect 2 -13 6 -9
<< pdcontact >>
rect -6 8 -2 12
rect 2 1 6 5
<< psubstratepcontact >>
rect -10 -20 -6 -16
<< nsubstratencontact >>
rect -10 8 -6 12
<< labels >>
rlabel metal1 7 10 7 10 6 Vdd!
rlabel metal1 7 -18 7 -18 7 Gnd!
rlabel polysilicon 0 -2 0 -2 1 A
rlabel metal1 5 -2 5 -2 7 F
<< end >>
